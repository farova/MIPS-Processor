`ifndef _control_vh_
`define _control_vh_

`define CNTRL_REG_SIZE 17

`define BR 0
`define JP 1
`define DMWE 2
`define RWE 3
`define RWD 4
`define RDST 5
`define ALUOP 6
`define ALUINB 7
`define JR 8
`define RA 9
`define BYTE 10
`define UBYTE 11
`define SRC1 12
`define SRC2 13
`define DEST 14
`define LOAD 15
`define STORE 16

`endif 