module Execute();

endmodule