`ifndef _control_vh_
`define _control_vh_

`define CNTRL_REG_SIZE 12

`define BR 0
`define JP 1
`define DMWE 2
`define RWE 3
`define RWD 4
`define RDST 5
`define ALUOP 6
`define ALUINB 7
`define JR 8
`define RA 9
`define BYTE 10
`define UBYTE 11

`endif 